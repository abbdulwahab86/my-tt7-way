module rom_S9(
    input wire [8:0] address,
    output reg [8:0] data
);

// Memory content initialization
reg [8:0] memory [511:0]; // 2^9 = 512 locations;memory[] = 9'dindexed from 0 to 511

// Initialize memory content with provided values
initial 
begin

memory[0] = 9'd167;
memory[1] = 9'd239;
memory[2] = 9'd161;
memory[3] = 9'd379;
memory[4] = 9'd391;
memory[5] = 9'd334;
memory[6] = 9'd9;
memory[7] = 9'd338;
memory[8] = 9'd38;
memory[9] = 9'd226;
memory[10] = 9'd48;
memory[11] = 9'd358;
memory[12] = 9'd452;
memory[13] = 9'd385;
memory[14] = 9'd90;
memory[15] = 9'd397;
memory[16] = 9'd183;
memory[17] = 9'd253;
memory[18] = 9'd147;
memory[19] = 9'd331;
memory[20] = 9'd415;
memory[21] = 9'd340;
memory[22] = 9'd51;
memory[23] = 9'd362;
memory[24] = 9'd306;
memory[25] = 9'd500;
memory[26] = 9'd262;
memory[27] = 9'd82;
memory[28] = 9'd216;
memory[29] = 9'd159;
memory[30] = 9'd356;
memory[31] = 9'd177;
memory[32] = 9'd175;
memory[33] = 9'd241;
memory[34] = 9'd489;
memory[35] = 9'd37;
memory[36] = 9'd206;
memory[37] = 9'd17;
memory[38] = 9'd0;
memory[39] = 9'd333;
memory[40] = 9'd44;
memory[41] = 9'd254;
memory[42] = 9'd378;
memory[43] = 9'd58;
memory[44] = 9'd143;
memory[45] = 9'd220;
memory[46] = 9'd81;
memory[47] = 9'd400;
memory[48] = 9'd95;
memory[49] = 9'd3;
memory[50] = 9'd315;
memory[51] = 9'd245;
memory[52] = 9'd54;
memory[53] = 9'd235;
memory[54] = 9'd218;
memory[55] = 9'd405;
memory[56] = 9'd472;
memory[57] = 9'd264;
memory[58] = 9'd172;
memory[59] = 9'd494;
memory[60] = 9'd371;
memory[61] = 9'd290;
memory[62] = 9'd399;
memory[63] = 9'd76;
memory[64] = 9'd165;
memory[65] = 9'd197;
memory[66] = 9'd395;
memory[67] = 9'd121;
memory[68] = 9'd257;
memory[69] = 9'd480;
memory[70] = 9'd423;
memory[71] = 9'd212;
memory[72] = 9'd240;
memory[73] = 9'd28;
memory[74] = 9'd462;
memory[75] = 9'd176;
memory[76] = 9'd406;
memory[77] = 9'd507;
memory[78] = 9'd288;
memory[79] = 9'd223;
memory[80] = 9'd501;
memory[81] = 9'd407;
memory[82] = 9'd249;
memory[83] = 9'd265;
memory[84] = 9'd89;
memory[85] = 9'd186;
memory[86] = 9'd221;
memory[87] = 9'd428;
memory[88] = 9'd164;
memory[89] = 9'd74;
memory[90] = 9'd440;
memory[91] = 9'd196;
memory[92] = 9'd458;
memory[93] = 9'd421;
memory[94] = 9'd350;
memory[95] = 9'd163;
memory[96] = 9'd232;
memory[97] = 9'd158;
memory[98] = 9'd134;
memory[99] = 9'd354;
memory[100] = 9'd13;
memory[101] = 9'd250;
memory[102] = 9'd491;
memory[103] = 9'd142;
memory[104] = 9'd191;
memory[105] = 9'd69;
memory[106] = 9'd193;
memory[107] = 9'd425;
memory[108] = 9'd152;
memory[109] = 9'd227;
memory[110] = 9'd366;
memory[111] = 9'd135;
memory[112] = 9'd344;
memory[113] = 9'd300;
memory[114] = 9'd276;
memory[115] = 9'd242;
memory[116] = 9'd437;
memory[117] = 9'd320;
memory[118] = 9'd113;
memory[119] = 9'd278;
memory[120] = 9'd11;
memory[121] = 9'd243;
memory[122] = 9'd87;
memory[123] = 9'd317;
memory[124] = 9'd36;
memory[125] = 9'd93;
memory[126] = 9'd496;
memory[127] = 9'd27;
memory[128] = 9'd487;
memory[129] = 9'd446;
memory[130] = 9'd482;
memory[131] = 9'd41;
memory[132] = 9'd68;
memory[133] = 9'd156;
memory[134] = 9'd457;
memory[135] = 9'd131;
memory[136] = 9'd326;
memory[137] = 9'd403;
memory[138] = 9'd339;
memory[139] = 9'd20;
memory[140] = 9'd39;
memory[141] = 9'd115;
memory[142] = 9'd442;
memory[143] = 9'd124;
memory[144] = 9'd475;
memory[145] = 9'd384;
memory[146] = 9'd508;
memory[147] = 9'd53;
memory[148] = 9'd112;
memory[149] = 9'd170;
memory[150] = 9'd479;
memory[151] = 9'd151;
memory[152] = 9'd126;
memory[153] = 9'd169;
memory[154] = 9'd73;
memory[155] = 9'd268;
memory[156] = 9'd279;
memory[157] = 9'd321;
memory[158] = 9'd168;
memory[159] = 9'd364;
memory[160] = 9'd363;
memory[161] = 9'd292;
memory[162] = 9'd46;
memory[163] = 9'd499;
memory[164] = 9'd393;
memory[165] = 9'd327;
memory[166] = 9'd324;
memory[167] = 9'd24;
memory[168] = 9'd456;
memory[169] = 9'd267;
memory[170] = 9'd157;
memory[171] = 9'd460;
memory[172] = 9'd488;
memory[173] = 9'd426;
memory[174] = 9'd309;
memory[175] = 9'd229;
memory[176] = 9'd439;
memory[177] = 9'd506;
memory[178] = 9'd208;
memory[179] = 9'd271;
memory[180] = 9'd349;
memory[181] = 9'd401;
memory[182] = 9'd434;
memory[183] = 9'd236;
memory[184] = 9'd16;
memory[185] = 9'd209;
memory[186] = 9'd359;
memory[187] = 9'd52;
memory[188] = 9'd56;
memory[189] = 9'd120;
memory[190] = 9'd199;
memory[191] = 9'd277;
memory[192] = 9'd465;
memory[193] = 9'd416;
memory[194] = 9'd252;
memory[195] = 9'd287;
memory[196] = 9'd246;
memory[197] = 9'd 6;
memory[198] = 9'd83;
memory[199] = 9'd305;
memory[200] = 9'd420;
memory[201] = 9'd345;
memory[202] = 9'd153;
memory[203] = 9'd502;
memory[204] = 9'd65;
memory[205] = 9'd61;
memory[206] = 9'd244;
memory[207] = 9'd282;
memory[208] = 9'd173;
memory[209] = 9'd222;
memory[210] = 9'd418;
memory[211] = 9'd67;
memory[212] = 9'd386;
memory[213] = 9'd368;
memory[214] = 9'd261;
memory[215] = 9'd101;
memory[216] = 9'd476;
memory[217] = 9'd291;
memory[218] = 9'd195;
memory[219] = 9'd430;
memory[220] = 9'd49;
memory[221] = 9'd79;
memory[222] = 9'd166;
memory[223] = 9'd330;
memory[224] = 9'd280;
memory[225] = 9'd383;
memory[226] = 9'd373;
memory[227] = 9'd128;
memory[228] = 9'd382;
memory[229] = 9'd408;
memory[230] = 9'd155;
memory[231] = 9'd495;
memory[232] = 9'd367;
memory[233] = 9'd388;
memory[234] = 9'd274;
memory[235] = 9'd107;
memory[236] = 9'd459;
memory[237] = 9'd417;
memory[238] = 9'd62;
memory[239] = 9'd454;
memory[240] = 9'd132;
memory[241] = 9'd225;
memory[242] = 9'd203;
memory[243] = 9'd316;
memory[244] = 9'd234;
memory[245] = 9'd14;
memory[246] = 9'd301;
memory[247] = 9'd91;
memory[248] = 9'd503;
memory[249] = 9'd286;
memory[250] = 9'd424;
memory[251] = 9'd211;
memory[252] = 9'd347;
memory[253] = 9'd307;
memory[254] = 9'd140;
memory[255] = 9'd374;
memory[256] = 9'd35;
memory[257] = 9'd103;
memory[258] = 9'd125;
memory[259] = 9'd427;
memory[260] = 9'd19;
memory[261] = 9'd214;
memory[262] = 9'd453;
memory[263] = 9'd146;
memory[264] = 9'd498;
memory[265] = 9'd314;
memory[266] = 9'd444;
memory[267] = 9'd230;
memory[268] = 9'd256;
memory[269] = 9'd329;
memory[270] = 9'd198;
memory[271] = 9'd285;
memory[272] = 9'd50;
memory[273] = 9'd116;
memory[274] = 9'd78;
memory[275] = 9'd410;
memory[276] = 9'd10;
memory[277] = 9'd205;
memory[278] = 9'd510;
memory[279] = 9'd171;
memory[280] = 9'd231;
memory[281] = 9'd45;
memory[282] = 9'd139;
memory[283] = 9'd467;
memory[284] = 9'd29;
memory[285] = 9'd86;
memory[286] = 9'd505;
memory[287] = 9'd32;
memory[288] = 9'd72;
memory[289] = 9'd26;
memory[290] = 9'd342;
memory[291] = 9'd150;
memory[292] = 9'd313;
memory[293] = 9'd490;
memory[294] = 9'd431;
memory[295] = 9'd238;
memory[296] = 9'd411;
memory[297] = 9'd325;
memory[298] = 9'd149;
memory[299] = 9'd473;
memory[300] = 9'd40;
memory[301] = 9'd119;
memory[302] = 9'd174;
memory[303] = 9'd355;
memory[304] = 9'd185;
memory[305] = 9'd233;
memory[306] = 9'd389;
memory[307] = 9'd71;
memory[308] = 9'd448;
memory[309] = 9'd273;
memory[310] = 9'd372;
memory[311] = 9'd55;
memory[312] = 9'd110;
memory[313] = 9'd178;
memory[314] = 9'd322;
memory[315] = 9'd12;
memory[316] = 9'd469;
memory[317] = 9'd392;
memory[318] = 9'd369;
memory[319] = 9'd190;
memory[320] = 9'd1;
memory[321] = 9'd109;
memory[322] = 9'd375;
memory[323] = 9'd137;
memory[324] = 9'd181;
memory[325] = 9'd88;
memory[326] = 9'd75;
memory[327] = 9'd308;
memory[328] = 9'd260;
memory[329] = 9'd484;
memory[330] = 9'd98;
memory[331] = 9'd272;
memory[332] = 9'd370;
memory[333] = 9'd275;
memory[334] = 9'd412;
memory[335] = 9'd111;
memory[336] = 9'd336;
memory[337] = 9'd318;
memory[338] = 9'd4;
memory[339] = 9'd504;
memory[340] = 9'd492;
memory[341] = 9'd259;
memory[342] = 9'd304;
memory[343] = 9'd77;
memory[344] = 9'd337;
memory[345] = 9'd435;
memory[346] = 9'd21;
memory[347] = 9'd357;
memory[348] = 9'd303;
memory[349] = 9'd332;
memory[350] = 9'd483;
memory[351] = 9'd18;
memory[352] = 9'd47;
memory[353] = 9'd85;
memory[354] = 9'd25;
memory[355] = 9'd497;
memory[356] = 9'd474;
memory[357] = 9'd289;
memory[358] = 9'd100;
memory[359] = 9'd269;
memory[360] = 9'd296;
memory[361] = 9'd478;
memory[362] = 9'd270;
memory[363] = 9'd106;
memory[364] = 9'd31;
memory[365] = 9'd104;
memory[366] = 9'd433;
memory[367] = 9'd84;
memory[368] = 9'd414;
memory[369] = 9'd486;
memory[370] = 9'd394;
memory[371] = 9'd96;
memory[372] = 9'd99;
memory[373] = 9'd154;
memory[374] = 9'd511;
memory[375] = 9'd148;
memory[376] = 9'd413;
memory[377] = 9'd361;
memory[378] = 9'd409;
memory[379] = 9'd255;
memory[380] = 9'd162;
memory[381] = 9'd215;
memory[382] = 9'd302;
memory[383] = 9'd201;
memory[384] = 9'd266;
memory[385] = 9'd351;
memory[386] = 9'd343;
memory[387] = 9'd144;
memory[388] = 9'd441;
memory[389] = 9'd365;
memory[390] = 9'd108;
memory[391] = 9'd298;
memory[392] = 9'd251;
memory[393] = 9'd34;
memory[394] = 9'd182;
memory[395] = 9'd509;
memory[396] = 9'd138;
memory[397] = 9'd210;
memory[398] = 9'd335;
memory[399] = 9'd133;
memory[400] = 9'd311;
memory[401] = 9'd352;
memory[402] = 9'd328;
memory[403] = 9'd141;
memory[404] = 9'd396;
memory[405] = 9'd346;
memory[406] = 9'd123;
memory[407] = 9'd319;
memory[408] = 9'd450;
memory[409] = 9'd281;
memory[410] = 9'd429;
memory[411] = 9'd228;
memory[412] = 9'd443;
memory[413] = 9'd481;
memory[414] = 9'd92;
memory[415] = 9'd404;
memory[416] = 9'd485;
memory[417] = 9'd422;
memory[418] = 9'd248;
memory[419] = 9'd297;
memory[420] = 9'd23;
memory[421] = 9'd213;
memory[422] = 9'd130;
memory[423] = 9'd466;
memory[424] = 9'd22;
memory[425] = 9'd217;
memory[426] = 9'd283;
memory[427] = 9'd70;
memory[428] = 9'd294;
memory[429] = 9'd360;
memory[430] = 9'd419;
memory[431] = 9'd127;
memory[432] = 9'd312;
memory[433] = 9'd377;
memory[434] = 9'd7;
memory[435] = 9'd468;
memory[436] = 9'd194;
memory[437] = 9'd2;
memory[438] = 9'd117;
memory[439] = 9'd295;
memory[440] = 9'd463;
memory[441] = 9'd258;
memory[442] = 9'd224;
memory[443] = 9'd447;
memory[444] = 9'd247;
memory[445] = 9'd187;
memory[446] = 9'd80;
memory[447] = 9'd398;
memory[448] = 9'd284;
memory[449] = 9'd353;
memory[450] = 9'd105;
memory[451] = 9'd390;
memory[452] = 9'd299;
memory[453] = 9'd471;
memory[454] = 9'd470;
memory[455] = 9'd184;
memory[456] = 9'd57;
memory[457] = 9'd200;
memory[458] = 9'd348;
memory[459] = 9'd63;
memory[460] = 9'd204;
memory[461] = 9'd188;
memory[462] = 9'd33;
memory[463] = 9'd451;
memory[464] = 9'd97;
memory[465] = 9'd30;
memory[466] = 9'd310;
memory[467] = 9'd219;
memory[468] = 9'd94;
memory[469] = 9'd160;
memory[470] = 9'd129;
memory[471] = 9'd493;
memory[472] = 9'd64;
memory[473] = 9'd179;
memory[474] = 9'd263;
memory[475] = 9'd102;
memory[476] = 9'd189;
memory[477] = 9'd207;
memory[478] = 9'd114;
memory[479] = 9'd402;
memory[480] = 9'd438;
memory[481] = 9'd477;
memory[482] = 9'd387;
memory[483] = 9'd122;
memory[484] = 9'd192;
memory[485] = 9'd42;
memory[486] = 9'd381;
memory[487] = 9'd5;
memory[488] = 9'd145;
memory[489] = 9'd118;
memory[490] = 9'd180;
memory[491] = 9'd449;
memory[492] = 9'd293;
memory[493] = 9'd323;
memory[494] = 9'd136;
memory[495] = 9'd380;
memory[496] = 9'd43;
memory[497] = 9'd66;
memory[498] = 9'd60;
memory[499] = 9'd455;
memory[500] = 9'd341;
memory[501] = 9'd445;
memory[502] = 9'd202;
memory[503] = 9'd432;
memory[504] = 9'd8;
memory[505] = 9'd237;
memory[506] = 9'd15;
memory[507] = 9'd376;
memory[508] = 9'd436;
memory[509] = 9'd464;
memory[510] = 9'd59;
memory[511] = 9'd461;
end
// Read operation
always @ (address)
    data <= memory[address];

endmodule